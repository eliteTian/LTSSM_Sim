`timescale 1ns/100ps
`include "define.v"
/* This project is aimed for understanding core LTSSM transition.
It's meant to be a digital only project, many core analog signals
are omitted or substituted by simulation construct. The core is
fully synthesizable and expandable and can be built into product IP
if expanded with enough features.*/
/*TS1 and TS2s are meant to be transmitted directly. The project is
two LTSSMs of same module talking to each other via TS1s. This process
simplifies the communication and eliminates the complexity of serdes
sim*/
/*TS1s are transmitted serially over the differential pair. The speed of
different gens are
Gen1: 2.5G/s    serial clock cycle and freq: 400ps 2.5GHz
Gen2: 5.0G/s    serial clock cycle and freq: 200ps 5.0GHz
Gen3: 8.0G/s    serial clock cycle and freq: 125ps 8.0GHz
Gen4: 16G/s     serial clock cycle and freq: 62.5ps 16.0GHz
Gen5: 32G/s     serial clock cycle and freq: 31.25ps 32.0GHz

Say system digital clock speed is 1GHz, the parallel TSs come in at a given
rate:
TS1: 16symbol = 128bit, Throughput = 128bitx1G = 128Gbps/per lane
assuming TS1s are sent back to back.
Gen1: 2.5Gx0.8(overhead) = 2Gbps. coming at 1 valid/ 128/2=64 cycles
Gen2: 5.0Gx0.8(overhead) = 4Gbps. coming at 1 valid/ 128/4=32 cycles
Gen3: 8.0Gx(128/130) = 8Gbps(neglecting encoding): coming at 1 valid/ 128/8=16 cycles
Gen4: 16.0Gx(128/130) = 16Gbps(neglecting encoding): coming at 1 valid/ 128/16=8 cycles
Gen5: 32.0Gx(128/130) = 32Gbps(neglecting encoding): coming at 1 valid/ 128/32=4 cycles

*/


module LTSSM(
    input            clk, //1GHz sys clock.
    input            rst,
    input            mode, //0:DSP, 1:USP
    //RX detect
    input            lane0_rx_det,
    input            lane1_rx_det,
    input            lane2_rx_det,
    input            lane3_rx_det,

    input            lane0_idle_break,
    input            lane1_idle_break,
    input            lane2_idle_break,
    input            lane3_idle_break,

    output           lane0_rx_det_seq_req,
    output           lane1_rx_det_seq_req,
    output           lane2_rx_det_seq_req,
    output           lane3_rx_det_seq_req,

    input            lane0_rx_det_seq_ack,
    input            lane1_rx_det_seq_ack,
    input            lane2_rx_det_seq_ack,
    input            lane3_rx_det_seq_ack,

    
    //TS1/s IF
    input[127:0]     lane0_ts_i,
    input            lane0_ts_i_vld,
    output[127:0]    lane0_ts_o,
    output           lane0_ts_o_vld,
    input[127:0]     lane1_ts_i,
    input            lane1_ts_i_vld,
    output[127:0]    lane1_ts_o,
    output           lane1_ts_o_vld,
    input[127:0]     lane2_ts_i,
    input            lane2_ts_i_vld,
    output[127:0]    lane2_ts_o,
    output           lane2_ts_o_vld,
    input[127:0]     lane3_ts_i,
    input            lane3_ts_i_vld,
    output[127:0]    lane3_ts_o,
    output           lane3_ts_o_vld,

    input            lane0_tx_fifo_full,
    input            lane1_tx_fifo_full,
    input            lane2_tx_fifo_full,
    input            lane3_tx_fifo_full,

    output[5:0]      curr_speed,
    output           linkup
);

wire[3:0]   w_elec_idle_brk     =   {lane3_idle_break,lane2_idle_break,lane1_idle_break,lane0_idle_break};
wire[3:0]   w_rx_det_seq_ack    =   {lane3_rx_det_seq_ack,lane2_rx_det_seq_ack,lane1_rx_det_seq_ack,lane0_rx_det_seq_ack};
wire[3:0]   w_rx_det_seq_req;
assign      {lane3_rx_det_seq_req,lane2_rx_det_seq_req,lane1_rx_det_seq_req,lane0_rx_det_seq_req} = w_rx_det_seq_req;

wire[3:0]   w_lanes_rx_det; 
assign      w_lanes_rx_det = {lane3_rx_det, lane2_rx_det, lane1_rx_det, lane0_rx_det} ;

wire[7:0]   w_ts_info;
wire        w_ts_update;

wire[3:0]   w_ts_update_ack_tx;
wire[3:0]   w_ts_update_ack_rx;

wire    lane0_sent_enough;
wire    lane1_sent_enough;
wire    lane2_sent_enough;
wire    lane3_sent_enough;

wire    lane0_tsa_p_a2c;
wire    lane1_tsa_p_a2c;
wire    lane2_tsa_p_a2c;
wire    lane3_tsa_p_a2c;

wire    lane0_tsa_p2c;
wire    lane1_tsa_p2c;
wire    lane2_tsa_p2c;
wire    lane3_tsa_p2c;

wire    lane3_tsa_c_lw_s2a;
wire    lane2_tsa_c_lw_s2a;
wire    lane1_tsa_c_lw_s2a;
wire    lane0_tsa_c_lw_s2a;
  

ts_gen ts_gen_u0(
   .clk                             (clk), //1GHz sys clock.
   .rst                             (rst),
   .ts_info                         (w_ts_info), //state:[7:4] sub_state[3:0]
   .ts_update                       (w_ts_update),
   .ts_update_ack                   (w_ts_update_ack_tx[0]),   
   .ts_stop                         (ts_stop),
   .lane_num                        (4'b0001),
   .mode                            (mode),
   .to_tsa_ts_sent_enough           (lane0_sent_enough),
   .ts_valid                        (lane0_ts_o_vld),
   .ts                              (lane0_ts_o),
   .ts_tx_fifo_full                 (lane0_tx_fifo_full)
);

tsa u_tsa_u0 (
    .clk                            (clk),                  // 1GHz system clock
    .rst                            (rst),
    .ts_info                        (w_ts_info),              // [7:4] state, [3:0] substate
    .ts_update                      (w_ts_update),
    .ts_update_ack                  (w_ts_update_ack_rx[0]),
    .ts_stop                        (ts_stop),
    .speed                          (speed),
    .lane_num                       (4'b0001),
    .mode                           (mode),
    .to_tsa_ts_sent_enough          (lane0_sent_enough), // controller info per substate
    .remote_ts_valid                (lane0_ts_i_vld), 
    .remote_ts                      (lane0_ts_i),            // 128-bit remote TS
    .tsa_p_a2c                      (lane0_tsa_p_a2c),
    .tsa_c_lw_s2a                   (lane0_tsa_c_lw_s2a),    
    .tsa_p2c                        (lane0_tsa_p2c)
    
);

ts_gen ts_gen_u1(
   .clk                             (clk), //1GHz sys clock.
   .rst                             (rst),
   .ts_info                         (w_ts_info), //state:[7:4] sub_state[3:0]
   .ts_update                       (w_ts_update),
   .ts_update_ack                   (w_ts_update_ack_tx[1]), 
   .ts_stop                         (ts_stop),    
   .lane_num                        (4'b0010), 
   .mode                            (mode),  
   .to_tsa_ts_sent_enough           (lane1_sent_enough),
   .ts_valid                        (lane1_ts_o_vld),
   .ts                              (lane1_ts_o),
   .ts_tx_fifo_full                 (lane1_tx_fifo_full)
);

tsa u_tsa_u1 (
    .clk                            (clk),                  // 1GHz system clock
    .rst                            (rst),
    .ts_info                        (w_ts_info),              // [7:4] state, [3:0] substate
    .ts_update                      (w_ts_update),
    .ts_update_ack                  (w_ts_update_ack_rx[1]),
    .ts_stop                        (ts_stop),
    .lane_num                       (4'b0010),
    .mode                           (mode),   
    .speed                          (speed),
    .to_tsa_ts_sent_enough          (lane1_sent_enough), // controller info per substate
    .remote_ts_valid                (lane1_ts_i_vld),
    .remote_ts                      (lane1_ts_i),            // 128-bit remote TS
    .tsa_p_a2c                      (lane1_tsa_p_a2c),
    .tsa_c_lw_s2a                   (lane1_tsa_c_lw_s2a),    
    .tsa_p2c                        (lane1_tsa_p2c)
    
);

ts_gen ts_gen_u2(
   .clk                             (clk), //1GHz sys clock.
   .rst                             (rst),
   .ts_info                         (w_ts_info), //state:[7:4] sub_state[3:0]
   .ts_update                       (w_ts_update),
   .ts_update_ack                   (w_ts_update_ack_tx[2]),
   .ts_stop                         (ts_stop),    
   .lane_num                        (4'b0100),   
   .mode                            (mode),
   .to_tsa_ts_sent_enough           (lane2_sent_enough),
   .ts_valid                        (lane2_ts_o_vld),
   .ts                              (lane2_ts_o),
   .ts_tx_fifo_full                 (lane2_tx_fifo_full)
);

tsa u_tsa_u2 (
    .clk                            (clk),                  // 1GHz system clock
    .rst                            (rst),
    .ts_info                        (w_ts_info),              // [7:4] state, [3:0] substate
    .ts_update                      (w_ts_update),
    .ts_update_ack                  (w_ts_update_ack_rx[2]),
    .ts_stop                        (ts_stop),
    .lane_num                       (4'b0100),
    .mode                           (mode),
    .speed                          (speed),
    .to_tsa_ts_sent_enough          (lane2_sent_enough), // controller info per substate
    .remote_ts_valid                (lane2_ts_i_vld),
    .remote_ts                      (lane2_ts_i),            // 128-bit remote TS
    .tsa_p_a2c                      (lane2_tsa_p_a2c),
    .tsa_c_lw_s2a                   (lane2_tsa_c_lw_s2a),    
    .tsa_p2c                        (lane2_tsa_p2c)
    
);

ts_gen ts_gen_u3(
   .clk                             (clk), //1GHz sys clock.
   .rst                             (rst),
   .ts_info                         (w_ts_info), //state:[7:4] sub_state[3:0]
   .ts_update                       (w_ts_update),
   .ts_update_ack                   (w_ts_update_ack_tx[3]),
   .ts_stop                         (ts_stop),
   .lane_num                        (4'b1000),
   .mode                            (mode),
   .to_tsa_ts_sent_enough           (lane3_sent_enough),
   .ts_valid                        (lane3_ts_o_vld),
   .ts                              (lane3_ts_o),
   .ts_tx_fifo_full                 (lane3_tx_fifo_full)
);

tsa u_tsa_u3 (
    .clk                            (clk),                  // 1GHz system clock
    .rst                            (rst),
    .ts_info                        (w_ts_info),              // [7:4] state, [3:0] substate
    .ts_update                      (w_ts_update),
    .ts_update_ack                  (w_ts_update_ack_rx[3]),
    .ts_stop                        (ts_stop),
    .speed                          (speed),
    .lane_num                       (4'b1000),
    .mode                           (mode),
    .to_tsa_ts_sent_enough          (lane3_sent_enough), // controller info per substate
    .remote_ts_valid                (lane3_ts_i_vld),
    .remote_ts                      (lane3_ts_i),            // 128-bit remote TS
    .tsa_p_a2c                      (lane3_tsa_p_a2c),
    .tsa_c_lw_s2a                   (lane3_tsa_c_lw_s2a),
    .tsa_p2c                        (lane3_tsa_p2c)
);

core_fsm core_fsm_u(
    .clk                            (clk), //1GHz sys clock.
    .rst                            (rst),
    .mode                           (mode),
    .elec_idle_break                (w_elec_idle_brk),
    .rx_det_seq_req                 (w_rx_det_seq_req),
    .rx_det_seq_ack                 (w_rx_det_seq_ack),
    .rx_det_valid                   (w_lanes_rx_det),

    .ts_info                        (w_ts_info), //state:[7:4] sub_state[3:0]
    .ts_update                      (w_ts_update),
    .ts_update_ack                  (w_ts_update_ack_tx&w_ts_update_ack_rx), //bitwise AND
    .ts_stop                        (w_ts_stop),
    
    .curr_speed                     (curr_speed),
    .tsa_p2c                        ({lane3_tsa_p2c , lane2_tsa_p2c , lane1_tsa_p2c , lane0_tsa_p2c}),
    .tsa_c_lw_s2a                   ({lane3_tsa_c_lw_s2a , lane2_tsa_c_lw_s2a , lane1_tsa_c_lw_s2a , lane0_tsa_c_lw_s2a}),
    .tsa_p_a2c                      ({lane3_tsa_p_a2c , lane2_tsa_p_a2c , lane1_tsa_p_a2c , lane0_tsa_p_a2c})
);

endmodule
    

