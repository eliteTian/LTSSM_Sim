`timescale 1ns/100ps
`include "define.v"
module core_fsm(
    input                    clk, //1GHz sys clock.
    input                    rst,
    input                    mode,
    //DETECT STATE
    input[`LANE_NUM-1:0]     elec_idle_break,
    output[`LANE_NUM-1:0]    rx_det_seq_req,
    input[`LANE_NUM-1:0]     rx_det_seq_ack,
    input[`LANE_NUM-1:0]     rx_det_valid,
    //POLL STATE
    output[7:0]              ts_info, //state:[7:4] sub_state[3:0]
    output                   ts_update,
    input[3:0]               ts_update_ack,
    output                   ts_stop,
    output[5:0]              curr_speed,
    //transition signals generated by ts analyzer
    input[`LANE_NUM-1:0]     tsa_p2c,    //polling to configuration
    input[`LANE_NUM-1:0]     tsa_p_a2c,   //polling active to polling configuration
    input[`LANE_NUM-1:0]     tsa_c_ws2wa,
    input[`LANE_NUM-1:0]     tsa_c_wa2nw


);

reg[31:0]                    cnt;
reg[31:0]                    timeout_val_reg, timeout_val_nxt;
reg                          cnt_start_reg, cnt_start_nxt;
reg                          pulse_set_reg, pulse_set_nxt;



reg[3:0]                     state_nxt, state_reg;
reg[1:0]                     detect_subst_nxt, detect_subst_reg;
reg[1:0]                     poll_subst_nxt, poll_subst_reg;
reg[3:0]                     cfg_subst_nxt, cfg_subst_reg;


reg[31:0]                    lane0_info_reg, lane1_info_reg, lane2_info_reg, lane3_info_reg;
reg[31:0]                    lane0_info_nxt, lane1_info_nxt, lane2_info_nxt, lane3_info_nxt;

reg[`LANE_NUM-1:0]           rx_det_seq_req_nxt, rx_det_seq_req_reg;
assign                       rx_det_seq_req = rx_det_seq_req_reg;

reg                          ts_update_nxt, ts_update_reg;
assign                       ts_update = ts_update_reg;

reg[7:0]                     ts_info_nxt, ts_info_reg;
assign                       ts_info = ts_info_reg;

//core LTSSM state transition.
always@(posedge clk) begin
    if(rst) begin
        state_reg <= `DETECT;
        detect_subst_reg <= `D_QUIET;
        poll_subst_reg <= `POLL_ACTIVE;
        cfg_subst_reg <= `CFG_LW_START;
    end else begin
        state_reg <= state_nxt;
        detect_subst_reg <= detect_subst_nxt;
        poll_subst_reg <= poll_subst_nxt;
        cfg_subst_reg <= cfg_subst_nxt;        
    end
end
//signals updating
always@(posedge clk) begin
    if(rst) begin
        pulse_set_reg <= `DETECT;
        cnt_start_reg <= 1'b0;
        timeout_val_reg <= 0;
        ts_info_reg <= 0;
        ts_update_reg <= 0;
        rx_det_seq_req_reg <= 0;
    end else begin
        pulse_set_reg <= pulse_set_nxt;
        cnt_start_reg <= cnt_start_nxt;
        timeout_val_reg <= timeout_val_nxt;
        ts_info_reg <= ts_info_nxt;
        ts_update_reg <= ts_update_nxt;
        rx_det_seq_req_reg <= rx_det_seq_req_nxt;
    end
end

/*state transition
Detect.quiet -> Detect.active : any lane has elec idle break. or 12ms timeout.
Detect.active -> Poll: 1.

*/
//
//down counter for generating timeout
always@(posedge clk) begin
    if(rst) begin
        cnt <= 32'hffffffff;
    end else begin
        if(cnt_start_reg) begin
            cnt <= timeout_val_reg;
        end /*else if(cnt_rst) begin
            cnt <= 0;
        end*/ else begin
            cnt <= cnt - 1;
        end
    end
end

wire timeout = ~|cnt & ~cnt_start_reg ;

always@* begin
    state_nxt = state_reg;
    detect_subst_nxt = detect_subst_reg;
    poll_subst_nxt = poll_subst_reg;
    cfg_subst_nxt = cfg_subst_reg;
    cnt_start_nxt = cnt_start_reg;
    timeout_val_nxt = timeout_val_reg;
    pulse_set_nxt = pulse_set_reg;
    ts_update_nxt = ts_update_reg;
    ts_info_nxt = ts_info_reg;
    rx_det_seq_req_nxt = rx_det_seq_req_reg;
    case(state_reg)
        `DETECT: begin
            case(detect_subst_reg)
                `D_QUIET: begin
                    if(~pulse_set_reg) begin //set counter, generate a single pulse to start counter
                        pulse_set_nxt = 1'b1;
                        cnt_start_nxt = 1'b1;
                        timeout_val_nxt = 'd12000000; //set as 12us to speed up sim;
                    end else begin
                        cnt_start_nxt = 1'b0;
                    end

                    if(|elec_idle_break || timeout) begin //@PCIe Gen5 Spec. 4.2.6.1.1 Detect.Quiet
                        detect_subst_nxt = `D_ACTIVE;
                        pulse_set_nxt = 1'b0;
                        rx_det_seq_req_nxt = 4'hF;
                    end
                end
                `D_ACTIVE: begin
                    if(~pulse_set_reg) begin //set counter, generate a single pulse to start counter
                        pulse_set_nxt = 1'b1;
                        cnt_start_nxt = 1'b1;
                        timeout_val_nxt = 'd12000; //set as 12us to speed up sim;
                    end else begin
                        cnt_start_nxt = 1'b0;
                    end

                    rx_det_seq_req_nxt = &rx_det_seq_ack ?  4'h0: rx_det_seq_req_reg ;

                    if(&rx_det_valid) begin //case 1, @PCIe Gen5 Spec. all lanes detect a valid receiver 4.2.6.1.2 Detect.Active
                        state_nxt = `POLL;
                        detect_subst_nxt = `D_QUIET;  
                        pulse_set_nxt = 1'b0;
                        rx_det_seq_req_nxt = 1'b0;
                    end

                    //if(~&rx_det_valid) begin //case 2, @PCIe Gen5 Spec. no lanes detect a valid receiver 4.2.6.1.2 Detect.Active
                    //    state_nxt = `DETECT;
                    //    detect_subst_nxt = `D_QUIET;  
                    //    pulse_set_nxt = 1'b0;
                    //    rx_det_seq_req_nxt = 1'b0;
                    //end // need to better monitor rx detect circuit, rx
                    //detect takes time and during this time, no state
                    //transition
                                            //cas3 3 to implement.
                    if(timeout) begin
                        detect_subst_nxt = `D_QUIET;
                    end
                end
            endcase
        end

        `POLL: begin
            case(poll_subst_reg)
                `POLL_ACTIVE: begin
                    if(~pulse_set_reg) begin //set timer, generate a single pulse to start counter
                        pulse_set_nxt = 1'b1;
                        cnt_start_nxt = 1'b1;
                        timeout_val_nxt = 'd24000; //set as 24us to speed up sim;
                        ts_info_nxt = {`POLL,`POLL_ACTIVE};//ts_info_nxt = {4'b0001,4'b0000};// ts_info_nxt = {`POLL,`POLL_ACTIVE};
                        ts_update_nxt = 1'b1;
                    end else begin
                        cnt_start_nxt = 1'b0;
                        ts_update_nxt = &ts_update_ack? 1'b0 :ts_update_reg ;
                    end

                    if(&tsa_p_a2c) begin
                        poll_subst_nxt = `POLL_CFG;
                        pulse_set_nxt = 1'b0;                        
                    end
                    if(timeout) begin
                        state_nxt = `DETECT;
                    end                    
                end
                `POLL_CFG: begin
                    if(~pulse_set_reg) begin //set timer, generate a single pulse to start counter
                        pulse_set_nxt = 1'b1;
                        cnt_start_nxt = 1'b1;
                        timeout_val_nxt = 'd24000; //set as 12us to speed up sim;
                        ts_info_nxt = {`POLL,`POLL_CFG};
                        ts_update_nxt = 1'b1;
                    end else begin
                        cnt_start_nxt = 1'b0;
                        ts_update_nxt = &ts_update_ack? 1'b0 :ts_update_reg ;
                    end

                    if(&tsa_p2c) begin
                        state_nxt = `CFG;
                        poll_subst_nxt = `POLL_ACTIVE;
                        pulse_set_nxt = 1'b0;
                    end
                    if(timeout) begin
                        state_nxt = `DETECT;
                    end
                end
            endcase
        end
        `CFG: begin
            case(cfg_subst_reg)
                `CFG_LW_START: begin
                    init_proc({`CFG,`CFG_LW_START},32'd24000);

                    if(&tsa_c_ws2wa) begin
                        cfg_subst_nxt = `CFG_LW_ACC;
                        pulse_set_nxt = 1'b0;
                    end
                    if(timeout) begin 
                        state_nxt = `DETECT;
                    end
                end

                `CFG_LW_ACC: begin
                    init_proc({`CFG,`CFG_LW_ACC},32'd24000);
                    if(&tsa_c_wa2nw) begin
                        cfg_subst_nxt = `CFG_LN_WAIT;
                        pulse_set_nxt = 1'b0;
                    end
                    if(timeout) begin 
                        state_nxt = `DETECT;
                    end
                end

                `CFG_LN_WAIT: begin
                    init_proc({`CFG,`CFG_LN_WAIT},32'd24000);


                    //if(&tsa_c_wa2na) begin
                    //    cfg_subst_nxt = `CFG_LN_ACC;
                    //    pulse_set_nxt = 1'b0;
                    //end
                    if(timeout) begin 
                        state_nxt = `DETECT;
                    end
                end




                //`CFG_COMPLETE: begin
                //    init_proc({`CFG,`CFG_LW_ACC},32'd24000);


                //    if(&tsa_c_wa2na) begin
                //        cfg_subst_nxt = `CFG_LN_WAIT;
                //        pulse_set_nxt = 1'b0;
                //    end
                //    if(timeout) begin 
                //        state_nxt = `DETECT;
                //    end
                //end






            endcase



        end
        
    endcase
end

assign curr_speed = `G1;

task init_proc;
input[7:0] ts_info;
input[31:0] timeout;
begin
    if(~pulse_set_reg) begin //set timer, generate a single pulse to start counter
        pulse_set_nxt = 1'b1;
        cnt_start_nxt = 1'b1;
        timeout_val_nxt = timeout; //set as 24us to speed up sim;
        ts_info_nxt = ts_info;
        ts_update_nxt = 1'b1;
    end else begin
        cnt_start_nxt = 1'b0;
        ts_update_nxt = &ts_update_ack? 1'b0 :ts_update_reg ;
    end
end
endtask

endmodule                  

